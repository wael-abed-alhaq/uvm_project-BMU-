`include "BMU_sequence_item.sv"
// `includBMUALU_random_SequeBMU
`include "BMU_interface.sv"

`include "BMU_reset_seq.sv"

`include "BMU_basic_operation_CSR_Bypass_Input_Data_seq.sv"
`include "csr_ren_in_apfields_not_zero_seq.sv"
`include "BMU_CSR_wr_data_ap_csr_imm_is_low_seq.sv"
`include "BMU_CSR_wr_data_ap_csr_imm_is_high_seq.sv"

`include "AND_operation_seq.sv"
`include "AND_operation_not_seq.sv"
`include "AND_operation_error_seq.sv"
`include "AND_operation_error2_seq.sv"
`include "OR_operation_seq.sv"
`include "OR_operation_not_seq.sv"
`include "OR_operation_error_seq.sv"
`include "OR_operation_error2_seq.sv"
`include "XOR_operation_seq.sv"
`include "XOR_operation_not_seq.sv"
`include "XOR_operation_error_seq.sv"
`include "XOR_operation_error2_seq.sv"

`include "sll_operation_basic_seq.sv"
`include "sll_operation_lower5_bits_in_bin_zero_seq.sv"
`include "sll_operation_lower5_bits_in_bin_one_seq.sv"
`include "srl_operation_basic_seq.sv"
`include "srl_operation_lower5_bits_in_bin_zero_seq.sv"
`include "srl_operation_lower5_bits_in_bin_one_seq.sv"
`include "sra_operation_basic_seq.sv"
`include "sra_operation_lower5_bits_in_bin_zero_seq.sv"
`include "sra_operation_lower5_bits_in_bin_one_seq.sv"
`include "rol_operation_basic_seq.sv"
`include "rol_operation_lower5_bits_in_bin_zero_seq.sv"
`include "rol_operation_lower5_bits_in_bin_one_seq.sv"
`include "ror_operation_basic_seq.sv"
`include "ror_operation_lower5_bits_in_bin_zero_seq.sv"
`include "ror_operation_lower5_bits_in_bin_one_seq.sv"
`include "bext_operation_basic_seq.sv"
`include "bext_operation_lower5_bits_in_bin_zero_seq.sv"
`include "bext_operation_lower5_bits_in_bin_one_seq.sv"
`include "binv_operation_basic_seq.sv"
`include "binv_operation_lower5_bits_in_bin_zero_seq.sv"
`include "binv_operation_lower5_bits_in_bin_one_seq.sv"
`include "sh1add_basic_seq.sv"
`include "sh1add_random_seq.sv"
`include "sh1add_error_seq.sv"
`include "sh2add_basic_seq.sv"
`include "sh2add_random_seq.sv"
`include "sh2add_error_seq.sv"
`include "sh3add_basic_seq.sv"
`include "sh3add_random_seq.sv"
`include "sh3add_error_seq.sv"

`include "subtract_seq.sv"
`include "subtract_error_seq.sv"
`include "ADD_seq.sv"
`include "ADD_overflow_seq.sv"

`include "set_on_less_than_seq.sv"
`include "clz_seq.sv"
`include "clz_input_zero_seq.sv"
`include "clz_input_most_significat_1_seq.sv"
`include "ctz_seq.sv"
`include "ctz_input_zero_seq.sv"
`include "ctz_input_least_significat_1_seq.sv"
`include "cpop_seq.sv"
`include "cpop_ain_zero_seq.sv"
`include "cpop_ain_ones_seq.sv"
`include "siext_b_seq.sv"
`include "siext_h_seq.sv"
`include "max_seq.sv"
`include "min_seq.sv"
`include "pack_seq.sv"
`include "packu_seq.sv"
`include "packh_seq.sv"
`include "grev_bin_24_seq.sv"
`include "grev_bin_not_24_seq.sv"
`include "gorc_basic_seq.sv"
`include "gorc_ain_zero_seq.sv"
`include "gorc_ain_ones_seq.sv"
`include "gorc_bin_not_7_seq.sv"
`include "gorc_ain_onebyte0_seq.sv"




`include "ref_model_1.sv"
// `include "BMU_add_sequence.sv"
// `include "BMU_sub_Sequence.sv"
// `includBMUALU_and_sequence.sv"
// `includBMUALU_or_sequence.sv"
// `includBMUALU_xor_sequence.sv"
// `includBMUALU_undefiend_opcode_sequence.sv"
// `includBMUALU_overflow_sequence.sv"
// `includBMUALU_underflow_Sequence.sv"
`include "BMU_sequencer.sv"
`include "BMU_driver.sv"
`include "BMU_monitor.sv"
`include "BMU_scoreboard.sv"
`include "BMU_subscriber.sv"
`include "BMU_agent.sv"
`include "BMU_enviroment.sv"
`include "BMU_base_test.sv"
`include "Control_Status_Reg_Oper_test.sv"
`include "Logic_operation_test.sv"
`include "BMU_shift_masking_operation_test.sv"
`include "BMU_Arithmetic_Operations_test.sv"
`include "Bit_Manipulation_test.sv"

